-- pragma translate_off
use std.textio.all;
-- pragma translate_on
package version is
  constant grlib_version : integer := 1021;
-- pragma translate_off
  constant grlib_date : string := "20090901";
-- pragma translate_on
  constant grlib_build : integer := 3848;
end;
